module alu (
    input wire [15:0] a,
    input wire [15:0] b,
    input wire [2:0] opcode,
    output wire [15:0] result,
    output wire zero,
    output wire carry
);
endmodule

