module counter (
    input wire clk,
    input wire reset,
    input wire enable,
    output wire [7:0] count
);
endmodule

