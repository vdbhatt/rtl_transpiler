module axi_crossbar (
    input wire aresetn,
    input wire [31:0] m0_awaddr,
    input wire [7:0] m0_awlen,
    input wire [2:0] m0_awsize,
    input wire [1:0] m0_awburst,
    input wire m0_awvalid,
    output wire m0_awready,
    input wire [63:0] m0_wdata,
    input wire [7:0] m0_wstrb,
    input wire m0_wlast,
    input wire m0_wvalid,
    output wire m0_wready,
    output wire [7:0] m0_bid,
    output wire [1:0] m0_bresp,
    output wire m0_bvalid,
    input wire m0_bready,
    input wire [7:0] m0_arid,
    input wire [31:0] m0_araddr,
    input wire [7:0] m0_arlen,
    input wire [2:0] m0_arsize,
    input wire [1:0] m0_arburst,
    input wire m0_arvalid,
    output wire m0_arready,
    output wire [7:0] m0_rid,
    output wire [63:0] m0_rdata,
    output wire [1:0] m0_rresp,
    output wire m0_rlast,
    output wire m0_rvalid,
    input wire m0_rready,
    output wire [31:0] s0_awaddr,
    output wire [7:0] s0_awlen,
    output wire [2:0] s0_awsize,
    output wire [1:0] s0_awburst,
    output wire s0_awvalid,
    input wire s0_awready,
    output wire [63:0] s0_wdata,
    output wire [7:0] s0_wstrb,
    output wire s0_wlast,
    output wire s0_wvalid,
    input wire s0_wready,
    input wire [7:0] s0_bid,
    input wire [1:0] s0_bresp,
    input wire s0_bvalid,
    output wire s0_bready,
    output wire [7:0] s0_arid,
    output wire [31:0] s0_araddr,
    output wire [7:0] s0_arlen,
    output wire [2:0] s0_arsize,
    output wire [1:0] s0_arburst,
    output wire s0_arvalid,
    input wire s0_arready,
    input wire [7:0] s0_rid,
    input wire [63:0] s0_rdata,
    input wire [1:0] s0_rresp,
    input wire s0_rlast,
    input wire s0_rvalid,
    output wire s0_rready
);
endmodule

